library verilog;
use verilog.vl_types.all;
entity LidarFrameView_vlg_tst is
    generic(
        CLK_PERIOD      : integer := 20
    );
end LidarFrameView_vlg_tst;
